module basic_or(input [4:0] b, input [4:0] c, output [8:0] a);

	assign a = b | c;

endmodule

