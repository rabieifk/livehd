
module basic_add (input [7:0] a, input [7:0] b,
  output [7:0] usum);

  assign usum =          a + b;
endmodule
