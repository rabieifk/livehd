
module basic_add2i (input [7:0] a, input [7:0] b, input [7:0] c,
  output [7:0] usum);

  assign usum =          a + b + c;
endmodule
