
module basic_sub (input [7:0] a, input [7:0] b,
output [7:0] usub);

  assign usub =          a - b;
endmodule
